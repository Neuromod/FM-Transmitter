module Loopback(rx, tx);
    input  wire rx;
    output wire tx;

    assign tx = rx;
endmodule
